module INTERPOLATION (    input               clk     ,    input               rst     ,    input   [  4:0]     frac_h  ,    input   [  4:0]     frac_w  ,    input   [  7:0]     d0      ,    input   [  7:0]     d1      ,    input   [  7:0]     d2      ,    input   [  7:0]     d3      ,    input               i_vld   ,    output  [  7:0]     o_d     ,    output              o_vld);reg     [ 12:0]     r_tmp0          ;reg     [  7:0]     r_tmp1          ;reg     [ 12:0]     r_tmp2          ;reg     [  7:0]     r_tmp3          ;reg     [  4:0]     r_frac_w        ;reg                 r_d1d0_plus     ;reg                 r_d3d2_plus     ;reg     [ 12:0]     r_tmp0_d0       ;reg     [ 15:0]     r_tmp1_d0       ;reg     [ 12:0]     r_tmp2_d0       ;reg     [ 15:0]     r_tmp3_d0       ;reg                 r_d1d0_plus_d0  ;reg                 r_d3d2_plus_d0  ;reg     [ 13:0]     r_d4            ;reg     [ 13:0]     r_d5            ;reg     [ 13:0]     r_d4_d0         ;reg     [ 13:0]     r_d5_d0         ;reg                 r_d5d4_plus     ;reg     [ 13:0]     r_d4_d1         ;reg     [ 16:0]     r_d5_d1         ;reg                 r_d5d4_plus_d0  ;reg     [ 13:0]     r_new_img       ;reg     [  5:0]     r_step_vld      ;wire                s_d1d0_plus     ;wire    [  7:0]     s_d1_d0         ;wire                s_d3d2_plus     ;wire    [  7:0]     s_d3_d2         ;wire                s_d5d4_plus     ;wire    [ 13:0]     s_d5_d4         ;always @ (posedge clk) begin    //step 0    r_tmp0          <= d0 << 5;    r_tmp1          <= s_d1_d0;    r_tmp2          <= d2 << 5;    r_tmp3          <= s_d3_d2;    r_frac_w        <= frac_w;    r_d1d0_plus     <= s_d1d0_plus;    r_d3d2_plus     <= s_d3d2_plus;    //step 1    r_tmp0_d0       <= r_tmp0;    r_tmp1_d0       <= r_tmp1 * r_frac_w;    r_tmp2_d0       <= r_tmp2;    r_tmp3_d0       <= r_tmp3 * r_frac_w;    r_d1d0_plus_d0  <= r_d1d0_plus;    r_d3d2_plus_d0  <= r_d3d2_plus;    //step 2    r_d4            <= r_d1d0_plus_d0 ? {3'd0,r_tmp0_d0} + r_tmp1_d0 : {3'd0,r_tmp0_d0} - r_tmp1_d0;    r_d5            <= r_d3d2_plus_d0 ? {3'd0,r_tmp2_d0} + r_tmp3_d0 : {3'd0,r_tmp2_d0} - r_tmp3_d0;    //step 3            r_d4_d0         <= r_d4;    r_d5_d0         <= s_d5_d4;    r_d5d4_plus     <= s_d5d4_plus;    //step 4    r_d4_d1         <= r_d4_d0;    r_d5_d1         <= r_d5_d0[13:5] * frac_h;     r_d5d4_plus_d0  <= r_d5d4_plus;    //step 5    r_new_img       <= r_d5d4_plus_d0 ? r_d4_d1 + r_d5_d1 : r_d4_d1 - r_d5_d1;        //step flag    if (rst) begin        r_step_vld  <= 6'd0;    end else begin        r_step_vld  <= {r_step_vld[4:0], i_vld};    endendassign s_d1d0_plus = (d1 > d0);assign s_d1_d0     = s_d1d0_plus ? d1 - d0 : d0 - d1;assign s_d3d2_plus = (d3 > d2);assign s_d3_d2     = s_d3d2_plus ? d3 - d2 : d2 - d3;  assign s_d5d4_plus = (r_d5 > r_d4);                        assign s_d5_d4     = s_d5d4_plus ? r_d5 - r_d4 : r_d4 - r_d5;  assign o_d      = r_new_img[12:5];assign o_vld    = r_step_vld[5];endmodule